LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY wrkCount IS
    	PORT 
    	(

    	    ALL_0, TOGGLE, OPTIMAL : IN STD_LOGIC;
    	    IS_7, OPT_Q2, OPT_Q2' : OUT STD_LOGIC

 
    	);
END wrkCount;